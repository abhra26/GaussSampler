module grom_x(
    input clk,
    input [31:0] ADDR,
    input [31:0] Din,
    input Enable,
    input [1:0] CNTRL,
    output [31:0] read_data,
    output status
);

parameter CNTRL_READ = 2'b01;
parameter CNTRL_WRITE = 2'b10;
parameter CNTRL_IDLE = 2'b00;

reg [31:0] mem [0:511];
reg [31:0] data_out;
reg stat;

assign read_data = data_out;
assign status = stat;

initial begin
    data_out <= 32'b0;
    stat <= 1'b0;
end

/*
initial 
    begin : init
        data_out <= 32'b0;
        stat <= 1'b0;
        mem[32'h0] = 32'b10000000000000000000000000000101;
        mem[32'h1] = 32'b00000000000000000000000000001000;
        mem[32'h2] = 32'b00000000000000000000000000000001;
        mem[32'h3] = 32'b10000000000000000000000000000111;
        mem[32'h4] = 32'b00000000000000000000000000000100;
        mem[32'h5] = 32'b10000000000000000000000000000001;
        mem[32'h6] = 32'b00000000000000000000000000001100;
        mem[32'h7] = 32'b00000000000000000000000000000001;
        mem[32'h8] = 32'b00000000000000000000000000000011;
        mem[32'h9] = 32'b10000000000000000000000000000011;
        mem[32'ha] = 32'b00000000000000000000000000001001;
        mem[32'hb] = 32'b00000000000000000000000000001001;
        mem[32'hc] = 32'b10000000000000000000000000001011;
        mem[32'hd] = 32'b00000000000000000000000000000101;
        mem[32'he] = 32'b10000000000000000000000000000100;
        mem[32'hf] = 32'b10000000000000000000000000000001;
        mem[32'h10] = 32'b00000000000000000000000000000100;
        mem[32'h11] = 32'b00000000000000000000000000000101;
        mem[32'h12] = 32'b00000000000000000000000000000011;
        mem[32'h13] = 32'b10000000000000000000000000000001;
        mem[32'h14] = 32'b00000000000000000000000000000001;
        mem[32'h15] = 32'b10000000000000000000000000000001;
        mem[32'h16] = 32'b00000000000000000000000000001000;
        mem[32'h17] = 32'b10000000000000000000000000000001;
        mem[32'h18] = 32'b10000000000000000000000000000010;
        mem[32'h19] = 32'b10000000000000000000000000000010;
        mem[32'h1a] = 32'b00000000000000000000000000000010;
        mem[32'h1b] = 32'b00000000000000000000000000000011;
        mem[32'h1c] = 32'b00000000000000000000000000000100;
        mem[32'h1d] = 32'b10000000000000000000000000000011;
        mem[32'h1e] = 32'b00000000000000000000000000000001;
        mem[32'h1f] = 32'b10000000000000000000000000001000;
        mem[32'h20] = 32'b10000000000000000000000000000110;
        mem[32'h21] = 32'b10000000000000000000000000000101;
        mem[32'h22] = 32'b00000000000000000000000000000101;
        mem[32'h23] = 32'b10000000000000000000000000001010;
        mem[32'h24] = 32'b00000000000000000000000000000111;
        mem[32'h25] = 32'b00000000000000000000000000001110;
        mem[32'h26] = 32'b10000000000000000000000000000100;
        mem[32'h27] = 32'b10000000000000000000000000000111;
        mem[32'h28] = 32'b00000000000000000000000000000001;
        mem[32'h29] = 32'b10000000000000000000000000000110;
        mem[32'h2a] = 32'b10000000000000000000000000000011;
        mem[32'h2b] = 32'b00000000000000000000000000001000;
        mem[32'h2c] = 32'b00000000000000000000000000000010;
        mem[32'h2d] = 32'b00000000000000000000000000001001;
        mem[32'h2e] = 32'b00000000000000000000000000000011;
        mem[32'h2f] = 32'b10000000000000000000000000000001;
        mem[32'h30] = 32'b10000000000000000000000000001000;
        mem[32'h31] = 32'b00000000000000000000000000000011;
        mem[32'h32] = 32'b10000000000000000000000000001000;
        mem[32'h33] = 32'b00000000000000000000000000000101;
        mem[32'h34] = 32'b10000000000000000000000000000101;
        mem[32'h35] = 32'b00000000000000000000000000000001;
        mem[32'h36] = 32'b10000000000000000000000000000001;
        mem[32'h37] = 32'b10000000000000000000000000001001;
        mem[32'h38] = 32'b00000000000000000000000000000100;
        mem[32'h39] = 32'b00000000000000000000000000000111;
        mem[32'h3a] = 32'b10000000000000000000000000001000;
        mem[32'h3b] = 32'b00000000000000000000000000001000;
        mem[32'h3c] = 32'b00000000000000000000000000000001;
        mem[32'h3d] = 32'b00000000000000000000000000000011;
        mem[32'h3e] = 32'b10000000000000000000000000001000;
        mem[32'h3f] = 32'b00000000000000000000000000000001;
        mem[32'h40] = 32'b00000000000000000000000000000001;
        mem[32'h41] = 32'b10000000000000000000000000000001;
        mem[32'h42] = 32'b00000000000000000000000000000010;
        mem[32'h43] = 32'b00000000000000000000000000000010;
        mem[32'h44] = 32'b00000000000000000000000000000011;
        mem[32'h45] = 32'b10000000000000000000000000000110;
        mem[32'h46] = 32'b00000000000000000000000000001000;
        mem[32'h47] = 32'b00000000000000000000000000000011;
        mem[32'h48] = 32'b10000000000000000000000000001000;
        mem[32'h49] = 32'b00000000000000000000000000000101;
        mem[32'h4a] = 32'b10000000000000000000000000000001;
        mem[32'h4b] = 32'b00000000000000000000000000000001;
        mem[32'h4c] = 32'b10000000000000000000000000000001;
        mem[32'h4d] = 32'b00000000000000000000000000000010;
        mem[32'h4e] = 32'b00000000000000000000000000000100;
        mem[32'h4f] = 32'b00000000000000000000000000000011;
        mem[32'h50] = 32'b00000000000000000000000000000011;
        mem[32'h51] = 32'b10000000000000000000000000000011;
        mem[32'h52] = 32'b10000000000000000000000000001000;
        mem[32'h53] = 32'b10000000000000000000000000000001;
        mem[32'h54] = 32'b10000000000000000000000000000010;
        mem[32'h55] = 32'b10000000000000000000000000000011;
        mem[32'h56] = 32'b00000000000000000000000000000011;
        mem[32'h57] = 32'b10000000000000000000000000000001;
        mem[32'h58] = 32'b10000000000000000000000000001001;
        mem[32'h59] = 32'b10000000000000000000000000001000;
        mem[32'h5a] = 32'b00000000000000000000000000000001;
        mem[32'h5b] = 32'b10000000000000000000000000000111;
        mem[32'h5c] = 32'b00000000000000000000000000001001;
        mem[32'h5d] = 32'b10000000000000000000000000000101;
        mem[32'h5e] = 32'b10000000000000000000000000000011;
        mem[32'h5f] = 32'b00000000000000000000000000001110;
        mem[32'h60] = 32'b10000000000000000000000000000010;
        mem[32'h61] = 32'b10000000000000000000000000000010;
        mem[32'h62] = 32'b10000000000000000000000000001000;
        mem[32'h63] = 32'b10000000000000000000000000001000;
        mem[32'h64] = 32'b10000000000000000000000000000010;
        mem[32'h65] = 32'b10000000000000000000000000000001;
        mem[32'h66] = 32'b10000000000000000000000000000010;
        mem[32'h67] = 32'b00000000000000000000000000000110;
        mem[32'h68] = 32'b00000000000000000000000000000001;
        mem[32'h69] = 32'b10000000000000000000000000000010;
        mem[32'h6a] = 32'b10000000000000000000000000000111;
        mem[32'h6b] = 32'b00000000000000000000000000000110;
        mem[32'h6c] = 32'b00000000000000000000000000000101;
        mem[32'h6d] = 32'b10000000000000000000000000000010;
        mem[32'h6e] = 32'b10000000000000000000000000000010;
        mem[32'h6f] = 32'b00000000000000000000000000000011;
        mem[32'h70] = 32'b10000000000000000000000000000111;
        mem[32'h71] = 32'b10000000000000000000000000001000;
        mem[32'h72] = 32'b00000000000000000000000000000110;
        mem[32'h73] = 32'b10000000000000000000000000001001;
        mem[32'h74] = 32'b00000000000000000000000000001000;
        mem[32'h75] = 32'b10000000000000000000000000000100;
        mem[32'h76] = 32'b00000000000000000000000000000011;
        mem[32'h77] = 32'b10000000000000000000000000000010;
        mem[32'h78] = 32'b00000000000000000000000000000111;
        mem[32'h79] = 32'b00000000000000000000000000000100;
        mem[32'h7a] = 32'b00000000000000000000000000000001;
        mem[32'h7b] = 32'b00000000000000000000000000000001;
        mem[32'h7c] = 32'b10000000000000000000000000001000;
        mem[32'h7d] = 32'b10000000000000000000000000000010;
        mem[32'h7e] = 32'b00000000000000000000000000000011;
        mem[32'h7f] = 32'b00000000000000000000000000001000;
        mem[32'h80] = 32'b00000000000000000000000000001101;
        mem[32'h81] = 32'b00000000000000000000000000000001;
        mem[32'h82] = 32'b00000000000000000000000000000101;
        mem[32'h83] = 32'b10000000000000000000000000000100;
        mem[32'h84] = 32'b10000000000000000000000000000111;
        mem[32'h85] = 32'b10000000000000000000000000000110;
        mem[32'h86] = 32'b00000000000000000000000000000101;
        mem[32'h87] = 32'b00000000000000000000000000000111;
        mem[32'h88] = 32'b00000000000000000000000000000101;
        mem[32'h89] = 32'b10000000000000000000000000000011;
        mem[32'h8a] = 32'b10000000000000000000000000000011;
        mem[32'h8b] = 32'b00000000000000000000000000000101;
        mem[32'h8c] = 32'b00000000000000000000000000000010;
        mem[32'h8d] = 32'b10000000000000000000000000000010;
        mem[32'h8e] = 32'b00000000000000000000000000000110;
        mem[32'h8f] = 32'b10000000000000000000000000000010;
        mem[32'h90] = 32'b00000000000000000000000000000010;
        mem[32'h91] = 32'b10000000000000000000000000000001;
        mem[32'h92] = 32'b10000000000000000000000000000101;
        mem[32'h93] = 32'b10000000000000000000000000001000;
        mem[32'h94] = 32'b10000000000000000000000000000100;
        mem[32'h95] = 32'b10000000000000000000000000000010;
        mem[32'h96] = 32'b00000000000000000000000000001000;
        mem[32'h97] = 32'b10000000000000000000000000000101;
        mem[32'h98] = 32'b10000000000000000000000000000011;
        mem[32'h99] = 32'b00000000000000000000000000000001;
        mem[32'h9a] = 32'b00000000000000000000000000000101;
        mem[32'h9b] = 32'b00000000000000000000000000000100;
        mem[32'h9c] = 32'b00000000000000000000000000001000;
        mem[32'h9d] = 32'b10000000000000000000000000000100;
        mem[32'h9e] = 32'b00000000000000000000000000001000;
        mem[32'h9f] = 32'b00000000000000000000000000000111;
        mem[32'ha0] = 32'b00000000000000000000000000000010;
        mem[32'ha1] = 32'b00000000000000000000000000000100;
        mem[32'ha2] = 32'b10000000000000000000000000000011;
        mem[32'ha3] = 32'b00000000000000000000000000000010;
        mem[32'ha4] = 32'b10000000000000000000000000000001;
        mem[32'ha5] = 32'b10000000000000000000000000000011;
        mem[32'ha6] = 32'b00000000000000000000000000000101;
        mem[32'ha7] = 32'b00000000000000000000000000000010;
        mem[32'ha8] = 32'b10000000000000000000000000000100;
        mem[32'ha9] = 32'b00000000000000000000000000000011;
        mem[32'haa] = 32'b00000000000000000000000000000001;
        mem[32'hab] = 32'b10000000000000000000000000000101;
        mem[32'hac] = 32'b00000000000000000000000000000011;
        mem[32'had] = 32'b00000000000000000000000000001000;
        mem[32'hae] = 32'b00000000000000000000000000000011;
        mem[32'haf] = 32'b10000000000000000000000000000001;
        mem[32'hb0] = 32'b00000000000000000000000000000001;
        mem[32'hb1] = 32'b10000000000000000000000000000001;
        mem[32'hb2] = 32'b10000000000000000000000000000001;
        mem[32'hb3] = 32'b00000000000000000000000000001000;
        mem[32'hb4] = 32'b10000000000000000000000000000011;
        mem[32'hb5] = 32'b00000000000000000000000000000100;
        mem[32'hb6] = 32'b00000000000000000000000000000001;
        mem[32'hb7] = 32'b10000000000000000000000000001001;
        mem[32'hb8] = 32'b00000000000000000000000000001001;
        mem[32'hb9] = 32'b00000000000000000000000000000110;
        mem[32'hba] = 32'b10000000000000000000000000000001;
        mem[32'hbb] = 32'b10000000000000000000000000000110;
        mem[32'hbc] = 32'b00000000000000000000000000000111;
        mem[32'hbd] = 32'b10000000000000000000000000000100;
        mem[32'hbe] = 32'b10000000000000000000000000000001;
        mem[32'hbf] = 32'b00000000000000000000000000001000;
        mem[32'hc0] = 32'b00000000000000000000000000000001;
        mem[32'hc1] = 32'b10000000000000000000000000000011;
        mem[32'hc2] = 32'b00000000000000000000000000000001;
        mem[32'hc3] = 32'b00000000000000000000000000000001;
        mem[32'hc4] = 32'b00000000000000000000000000000100;
        mem[32'hc5] = 32'b10000000000000000000000000000001;
        mem[32'hc6] = 32'b10000000000000000000000000000001;
        mem[32'hc7] = 32'b10000000000000000000000000001000;
        mem[32'hc8] = 32'b10000000000000000000000000000110;
        mem[32'hc9] = 32'b10000000000000000000000000000110;
        mem[32'hca] = 32'b10000000000000000000000000001011;
        mem[32'hcb] = 32'b10000000000000000000000000001011;
        mem[32'hcc] = 32'b10000000000000000000000000000101;
        mem[32'hcd] = 32'b10000000000000000000000000000110;
        mem[32'hce] = 32'b00000000000000000000000000000010;
        mem[32'hcf] = 32'b00000000000000000000000000000101;
        mem[32'hd0] = 32'b10000000000000000000000000000101;
        mem[32'hd1] = 32'b00000000000000000000000000000001;
        mem[32'hd2] = 32'b00000000000000000000000000000101;
        mem[32'hd3] = 32'b00000000000000000000000000000010;
        mem[32'hd4] = 32'b10000000000000000000000000000011;
        mem[32'hd5] = 32'b10000000000000000000000000000111;
        mem[32'hd6] = 32'b00000000000000000000000000001000;
        mem[32'hd7] = 32'b00000000000000000000000000001001;
        mem[32'hd8] = 32'b10000000000000000000000000000001;
        mem[32'hd9] = 32'b10000000000000000000000000000001;
        mem[32'hda] = 32'b00000000000000000000000000000011;
        mem[32'hdb] = 32'b10000000000000000000000000000011;
        mem[32'hdc] = 32'b10000000000000000000000000000001;
        mem[32'hdd] = 32'b10000000000000000000000000000001;
        mem[32'hde] = 32'b00000000000000000000000000000100;
        mem[32'hdf] = 32'b10000000000000000000000000001001;
        mem[32'he0] = 32'b10000000000000000000000000001101;
        mem[32'he1] = 32'b10000000000000000000000000000001;
        mem[32'he2] = 32'b10000000000000000000000000001000;
        mem[32'he3] = 32'b10000000000000000000000000000100;
        mem[32'he4] = 32'b10000000000000000000000000000110;
        mem[32'he5] = 32'b00000000000000000000000000000001;
        mem[32'he6] = 32'b10000000000000000000000000000010;
        mem[32'he7] = 32'b00000000000000000000000000000001;
        mem[32'he8] = 32'b10000000000000000000000000000001;
        mem[32'he9] = 32'b10000000000000000000000000000001;
        mem[32'hea] = 32'b00000000000000000000000000001000;
        mem[32'heb] = 32'b00000000000000000000000000001001;
        mem[32'hec] = 32'b10000000000000000000000000000011;
        mem[32'hed] = 32'b00000000000000000000000000000010;
        mem[32'hee] = 32'b00000000000000000000000000000010;
        mem[32'hef] = 32'b00000000000000000000000000001000;
        mem[32'hf0] = 32'b00000000000000000000000000000010;
        mem[32'hf1] = 32'b00000000000000000000000000000010;
        mem[32'hf2] = 32'b00000000000000000000000000001000;
        mem[32'hf3] = 32'b10000000000000000000000000000010;
        mem[32'hf4] = 32'b10000000000000000000000000000011;
        mem[32'hf5] = 32'b00000000000000000000000000001000;
        mem[32'hf6] = 32'b00000000000000000000000000000101;
        mem[32'hf7] = 32'b00000000000000000000000000000001;
        mem[32'hf8] = 32'b10000000000000000000000000000001;
        mem[32'hf9] = 32'b10000000000000000000000000000100;
        mem[32'hfa] = 32'b10000000000000000000000000000111;
        mem[32'hfb] = 32'b00000000000000000000000000001011;
        mem[32'hfc] = 32'b10000000000000000000000000000011;
        mem[32'hfd] = 32'b00000000000000000000000000001011;
        mem[32'hfe] = 32'b10000000000000000000000000001001;
        mem[32'hff] = 32'b00000000000000000000000000000100;
        mem[32'h100] = 32'b00000000000000000000000000000001;
        mem[32'h101] = 32'b00000000000000000000000000000001;
        mem[32'h102] = 32'b00000000000000000000000000000001;
        mem[32'h103] = 32'b10000000000000000000000000000010;
        mem[32'h104] = 32'b10000000000000000000000000000101;
        mem[32'h105] = 32'b00000000000000000000000000000001;
        mem[32'h106] = 32'b00000000000000000000000000000001;
        mem[32'h107] = 32'b00000000000000000000000000000001;
        mem[32'h108] = 32'b10000000000000000000000000000001;
        mem[32'h109] = 32'b10000000000000000000000000001010;
        mem[32'h10a] = 32'b10000000000000000000000000000100;
        mem[32'h10b] = 32'b10000000000000000000000000000111;
        mem[32'h10c] = 32'b00000000000000000000000000000001;
        mem[32'h10d] = 32'b10000000000000000000000000001000;
        mem[32'h10e] = 32'b10000000000000000000000000001011;
        mem[32'h10f] = 32'b10000000000000000000000000001100;
        mem[32'h110] = 32'b10000000000000000000000000000010;
        mem[32'h111] = 32'b00000000000000000000000000000011;
        mem[32'h112] = 32'b00000000000000000000000000000011;
        mem[32'h113] = 32'b00000000000000000000000000000111;
        mem[32'h114] = 32'b10000000000000000000000000001001;
        mem[32'h115] = 32'b00000000000000000000000000000011;
        mem[32'h116] = 32'b10000000000000000000000000000010;
        mem[32'h117] = 32'b10000000000000000000000000000011;
        mem[32'h118] = 32'b10000000000000000000000000000111;
        mem[32'h119] = 32'b00000000000000000000000000000011;
        mem[32'h11a] = 32'b00000000000000000000000000000010;
        mem[32'h11b] = 32'b10000000000000000000000000000001;
        mem[32'h11c] = 32'b10000000000000000000000000000101;
        mem[32'h11d] = 32'b10000000000000000000000000001001;
        mem[32'h11e] = 32'b10000000000000000000000000000010;
        mem[32'h11f] = 32'b00000000000000000000000000000011;
        mem[32'h120] = 32'b10000000000000000000000000000011;
        mem[32'h121] = 32'b10000000000000000000000000000010;
        mem[32'h122] = 32'b00000000000000000000000000000010;
        mem[32'h123] = 32'b10000000000000000000000000000011;
        mem[32'h124] = 32'b10000000000000000000000000000101;
        mem[32'h125] = 32'b00000000000000000000000000001100;
        mem[32'h126] = 32'b10000000000000000000000000000010;
        mem[32'h127] = 32'b10000000000000000000000000000001;
        mem[32'h128] = 32'b10000000000000000000000000000001;
        mem[32'h129] = 32'b10000000000000000000000000000100;
        mem[32'h12a] = 32'b10000000000000000000000000000100;
        mem[32'h12b] = 32'b10000000000000000000000000000001;
        mem[32'h12c] = 32'b10000000000000000000000000000010;
        mem[32'h12d] = 32'b00000000000000000000000000000001;
        mem[32'h12e] = 32'b00000000000000000000000000000001;
        mem[32'h12f] = 32'b00000000000000000000000000001101;
        mem[32'h130] = 32'b00000000000000000000000000000100;
        mem[32'h131] = 32'b10000000000000000000000000000001;
        mem[32'h132] = 32'b10000000000000000000000000000011;
        mem[32'h133] = 32'b00000000000000000000000000000010;
        mem[32'h134] = 32'b10000000000000000000000000000110;
        mem[32'h135] = 32'b00000000000000000000000000001000;
        mem[32'h136] = 32'b00000000000000000000000000001001;
        mem[32'h137] = 32'b10000000000000000000000000000101;
        mem[32'h138] = 32'b10000000000000000000000000000001;
        mem[32'h139] = 32'b00000000000000000000000000000011;
        mem[32'h13a] = 32'b10000000000000000000000000000101;
        mem[32'h13b] = 32'b10000000000000000000000000000101;
        mem[32'h13c] = 32'b00000000000000000000000000000001;
        mem[32'h13d] = 32'b00000000000000000000000000000111;
        mem[32'h13e] = 32'b00000000000000000000000000000110;
        mem[32'h13f] = 32'b10000000000000000000000000000111;
        mem[32'h140] = 32'b00000000000000000000000000000011;
        mem[32'h141] = 32'b10000000000000000000000000000010;
        mem[32'h142] = 32'b10000000000000000000000000000101;
        mem[32'h143] = 32'b10000000000000000000000000000110;
        mem[32'h144] = 32'b10000000000000000000000000000001;
        mem[32'h145] = 32'b00000000000000000000000000000110;
        mem[32'h146] = 32'b00000000000000000000000000000010;
        mem[32'h147] = 32'b00000000000000000000000000001000;
        mem[32'h148] = 32'b00000000000000000000000000000001;
        mem[32'h149] = 32'b10000000000000000000000000000100;
        mem[32'h14a] = 32'b00000000000000000000000000000110;
        mem[32'h14b] = 32'b00000000000000000000000000000111;
        mem[32'h14c] = 32'b00000000000000000000000000000010;
        mem[32'h14d] = 32'b10000000000000000000000000000101;
        mem[32'h14e] = 32'b10000000000000000000000000000111;
        mem[32'h14f] = 32'b00000000000000000000000000001011;
        mem[32'h150] = 32'b00000000000000000000000000000100;
        mem[32'h151] = 32'b10000000000000000000000000000110;
        mem[32'h152] = 32'b00000000000000000000000000000111;
        mem[32'h153] = 32'b00000000000000000000000000000011;
        mem[32'h154] = 32'b00000000000000000000000000000101;
        mem[32'h155] = 32'b10000000000000000000000000000001;
        mem[32'h156] = 32'b10000000000000000000000000000011;
        mem[32'h157] = 32'b10000000000000000000000000001001;
        mem[32'h158] = 32'b00000000000000000000000000000100;
        mem[32'h159] = 32'b10000000000000000000000000000001;
        mem[32'h15a] = 32'b00000000000000000000000000000111;
        mem[32'h15b] = 32'b00000000000000000000000000001011;
        mem[32'h15c] = 32'b00000000000000000000000000001000;
        mem[32'h15d] = 32'b10000000000000000000000000000011;
        mem[32'h15e] = 32'b10000000000000000000000000000110;
        mem[32'h15f] = 32'b00000000000000000000000000000100;
        mem[32'h160] = 32'b00000000000000000000000000001110;
        mem[32'h161] = 32'b00000000000000000000000000000010;
        mem[32'h162] = 32'b00000000000000000000000000001010;
        mem[32'h163] = 32'b10000000000000000000000000000001;
        mem[32'h164] = 32'b10000000000000000000000000000010;
        mem[32'h165] = 32'b10000000000000000000000000000001;
        mem[32'h166] = 32'b10000000000000000000000000000010;
        mem[32'h167] = 32'b00000000000000000000000000000110;
        mem[32'h168] = 32'b10000000000000000000000000000011;
        mem[32'h169] = 32'b00000000000000000000000000000111;
        mem[32'h16a] = 32'b10000000000000000000000000000011;
        mem[32'h16b] = 32'b00000000000000000000000000001010;
        mem[32'h16c] = 32'b10000000000000000000000000001000;
        mem[32'h16d] = 32'b10000000000000000000000000001001;
        mem[32'h16e] = 32'b00000000000000000000000000000101;
        mem[32'h16f] = 32'b10000000000000000000000000000001;
        mem[32'h170] = 32'b10000000000000000000000000000011;
        mem[32'h171] = 32'b00000000000000000000000000000001;
        mem[32'h172] = 32'b00000000000000000000000000000100;
        mem[32'h173] = 32'b00000000000000000000000000001001;
        mem[32'h174] = 32'b10000000000000000000000000000011;
        mem[32'h175] = 32'b10000000000000000000000000000010;
        mem[32'h176] = 32'b10000000000000000000000000000011;
        mem[32'h177] = 32'b10000000000000000000000000000010;
        mem[32'h178] = 32'b00000000000000000000000000000100;
        mem[32'h179] = 32'b10000000000000000000000000000010;
        mem[32'h17a] = 32'b00000000000000000000000000001001;
        mem[32'h17b] = 32'b10000000000000000000000000000111;
        mem[32'h17c] = 32'b00000000000000000000000000001011;
        mem[32'h17d] = 32'b00000000000000000000000000001000;
        mem[32'h17e] = 32'b00000000000000000000000000000001;
        mem[32'h17f] = 32'b00000000000000000000000000000011;
        mem[32'h180] = 32'b10000000000000000000000000001000;
        mem[32'h181] = 32'b10000000000000000000000000000001;
        mem[32'h182] = 32'b00000000000000000000000000000111;
        mem[32'h183] = 32'b10000000000000000000000000000100;
        mem[32'h184] = 32'b10000000000000000000000000000010;
        mem[32'h185] = 32'b00000000000000000000000000000010;
        mem[32'h186] = 32'b00000000000000000000000000000010;
        mem[32'h187] = 32'b10000000000000000000000000000001;
        mem[32'h188] = 32'b00000000000000000000000000000001;
        mem[32'h189] = 32'b10000000000000000000000000000001;
        mem[32'h18a] = 32'b00000000000000000000000000001000;
        mem[32'h18b] = 32'b10000000000000000000000000000111;
        mem[32'h18c] = 32'b10000000000000000000000000000001;
        mem[32'h18d] = 32'b00000000000000000000000000000110;
        mem[32'h18e] = 32'b10000000000000000000000000000001;
        mem[32'h18f] = 32'b00000000000000000000000000000001;
        mem[32'h190] = 32'b00000000000000000000000000000110;
        mem[32'h191] = 32'b10000000000000000000000000001000;
        mem[32'h192] = 32'b10000000000000000000000000001001;
        mem[32'h193] = 32'b10000000000000000000000000000110;
        mem[32'h194] = 32'b00000000000000000000000000000001;
        mem[32'h195] = 32'b00000000000000000000000000000001;
        mem[32'h196] = 32'b00000000000000000000000000001010;
        mem[32'h197] = 32'b10000000000000000000000000000100;
        mem[32'h198] = 32'b10000000000000000000000000000010;
        mem[32'h199] = 32'b00000000000000000000000000000011;
        mem[32'h19a] = 32'b10000000000000000000000000000100;
        mem[32'h19b] = 32'b00000000000000000000000000001001;
        mem[32'h19c] = 32'b00000000000000000000000000000010;
        mem[32'h19d] = 32'b00000000000000000000000000000001;
        mem[32'h19e] = 32'b10000000000000000000000000000100;
        mem[32'h19f] = 32'b00000000000000000000000000000001;
        mem[32'h1a0] = 32'b00000000000000000000000000001000;
        mem[32'h1a1] = 32'b00000000000000000000000000000001;
        mem[32'h1a2] = 32'b00000000000000000000000000000001;
        mem[32'h1a3] = 32'b10000000000000000000000000000111;
        mem[32'h1a4] = 32'b00000000000000000000000000000001;
        mem[32'h1a5] = 32'b00000000000000000000000000000111;
        mem[32'h1a6] = 32'b00000000000000000000000000000010;
        mem[32'h1a7] = 32'b00000000000000000000000000000010;
        mem[32'h1a8] = 32'b10000000000000000000000000001000;
        mem[32'h1a9] = 32'b10000000000000000000000000000001;
        mem[32'h1aa] = 32'b00000000000000000000000000000110;
        mem[32'h1ab] = 32'b00000000000000000000000000000010;
        mem[32'h1ac] = 32'b00000000000000000000000000000001;
        mem[32'h1ad] = 32'b10000000000000000000000000000001;
        mem[32'h1ae] = 32'b00000000000000000000000000000100;
        mem[32'h1af] = 32'b00000000000000000000000000000011;
        mem[32'h1b0] = 32'b10000000000000000000000000001011;
        mem[32'h1b1] = 32'b10000000000000000000000000000001;
        mem[32'h1b2] = 32'b10000000000000000000000000000001;
        mem[32'h1b3] = 32'b10000000000000000000000000000111;
        mem[32'h1b4] = 32'b00000000000000000000000000000110;
        mem[32'h1b5] = 32'b10000000000000000000000000000001;
        mem[32'h1b6] = 32'b00000000000000000000000000000010;
        mem[32'h1b7] = 32'b00000000000000000000000000000101;
        mem[32'h1b8] = 32'b10000000000000000000000000000101;
        mem[32'h1b9] = 32'b00000000000000000000000000000101;
        mem[32'h1ba] = 32'b00000000000000000000000000000001;
        mem[32'h1bb] = 32'b00000000000000000000000000000111;
        mem[32'h1bc] = 32'b00000000000000000000000000000001;
        mem[32'h1bd] = 32'b10000000000000000000000000000110;
        mem[32'h1be] = 32'b00000000000000000000000000000001;
        mem[32'h1bf] = 32'b00000000000000000000000000000001;
        mem[32'h1c0] = 32'b10000000000000000000000000001000;
        mem[32'h1c1] = 32'b00000000000000000000000000000100;
        mem[32'h1c2] = 32'b00000000000000000000000000000100;
        mem[32'h1c3] = 32'b00000000000000000000000000000001;
        mem[32'h1c4] = 32'b10000000000000000000000000000001;
        mem[32'h1c5] = 32'b10000000000000000000000000000010;
        mem[32'h1c6] = 32'b10000000000000000000000000000011;
        mem[32'h1c7] = 32'b10000000000000000000000000000001;
        mem[32'h1c8] = 32'b10000000000000000000000000000011;
        mem[32'h1c9] = 32'b00000000000000000000000000000010;
        mem[32'h1ca] = 32'b00000000000000000000000000000010;
        mem[32'h1cb] = 32'b00000000000000000000000000000111;
        mem[32'h1cc] = 32'b00000000000000000000000000000010;
        mem[32'h1cd] = 32'b00000000000000000000000000001000;
        mem[32'h1ce] = 32'b10000000000000000000000000001001;
        mem[32'h1cf] = 32'b10000000000000000000000000000001;
        mem[32'h1d0] = 32'b00000000000000000000000000000010;
        mem[32'h1d1] = 32'b10000000000000000000000000000111;
        mem[32'h1d2] = 32'b10000000000000000000000000001110;
        mem[32'h1d3] = 32'b00000000000000000000000000001001;
        mem[32'h1d4] = 32'b10000000000000000000000000000010;
        mem[32'h1d5] = 32'b00000000000000000000000000000001;
        mem[32'h1d6] = 32'b00000000000000000000000000000110;
        mem[32'h1d7] = 32'b00000000000000000000000000000001;
        mem[32'h1d8] = 32'b00000000000000000000000000001001;
        mem[32'h1d9] = 32'b10000000000000000000000000000011;
        mem[32'h1da] = 32'b00000000000000000000000000000001;
        mem[32'h1db] = 32'b00000000000000000000000000000111;
        mem[32'h1dc] = 32'b00000000000000000000000000000011;
        mem[32'h1dd] = 32'b00000000000000000000000000000010;
        mem[32'h1de] = 32'b10000000000000000000000000000001;
        mem[32'h1df] = 32'b00000000000000000000000000000010;
        mem[32'h1e0] = 32'b00000000000000000000000000000110;
        mem[32'h1e1] = 32'b00000000000000000000000000000011;
        mem[32'h1e2] = 32'b10000000000000000000000000000001;
        mem[32'h1e3] = 32'b00000000000000000000000000001000;
        mem[32'h1e4] = 32'b00000000000000000000000000000010;
        mem[32'h1e5] = 32'b10000000000000000000000000001100;
        mem[32'h1e6] = 32'b10000000000000000000000000000100;
        mem[32'h1e7] = 32'b00000000000000000000000000000001;
        mem[32'h1e8] = 32'b10000000000000000000000000000101;
        mem[32'h1e9] = 32'b00000000000000000000000000000001;
        mem[32'h1ea] = 32'b00000000000000000000000000000011;
        mem[32'h1eb] = 32'b10000000000000000000000000001000;
        mem[32'h1ec] = 32'b10000000000000000000000000001001;
        mem[32'h1ed] = 32'b10000000000000000000000000000010;
        mem[32'h1ee] = 32'b10000000000000000000000000000011;
        mem[32'h1ef] = 32'b10000000000000000000000000001000;
        mem[32'h1f0] = 32'b00000000000000000000000000000010;
        mem[32'h1f1] = 32'b10000000000000000000000000000001;
        mem[32'h1f2] = 32'b00000000000000000000000000000011;
        mem[32'h1f3] = 32'b10000000000000000000000000000100;
        mem[32'h1f4] = 32'b10000000000000000000000000001000;
        mem[32'h1f5] = 32'b10000000000000000000000000001101;
        mem[32'h1f6] = 32'b10000000000000000000000000001000;
        mem[32'h1f7] = 32'b10000000000000000000000000000001;
        mem[32'h1f8] = 32'b10000000000000000000000000000100;
        mem[32'h1f9] = 32'b10000000000000000000000000000010;
        mem[32'h1fa] = 32'b00000000000000000000000000000001;
        mem[32'h1fb] = 32'b10000000000000000000000000001000;
        mem[32'h1fc] = 32'b10000000000000000000000000000010;
        mem[32'h1fd] = 32'b10000000000000000000000000001010;
        mem[32'h1fe] = 32'b10000000000000000000000000001110;
        mem[32'h1ff] = 32'b10000000000000000000000000001110;
               

    end
    
*/
    
always @(posedge clk) begin
    case (CNTRL)
        CNTRL_WRITE: 
            begin
                if (Enable) begin
                    mem[ADDR] <= Din;
                    stat <= 1'b1;
                end
            end
        CNTRL_READ:
            begin
                if (Enable) begin
                    data_out <=mem[ADDR];
                    stat <= 1'b1;
                end
            end
        CNTRL_IDLE:
            begin
                data_out <= 32'b0;
                stat <= 1'b0;
            end
    endcase
end

endmodule